<?xml version="1.0" encoding="UTF-8"?>
<Batch version="1.0"><TaskList><Task type="ResizeTask" enabled="True"><Width units="0">800</Width><Height units="0">300</Height><DPI>150</DPI><Filter>9</Filter><UseProportions>True</UseProportions></Task><Task type="SelAddTask" enabled="True"><Left units="0" base_point="0">966</Left><Right units="0" base_point="2">-557</Right><Top units="0" base_point="0">0</Top><Bottom units="0" base_point="2">0</Bottom><RoundWidth units="1">5</RoundWidth><RoundHeight units="1">5</RoundHeight><Type>0</Type><Operation>0</Operation><Intensity>255</Intensity></Task><Task type="WatermarkTask" enabled="True"><FileName><![CDATA[C:\Program Files (x86)\ImBatch\Graphics\Logo1.png]]></FileName><Transparency>100</Transparency><Mode>0</Mode><ResampleFilter>0</ResampleFilter><Operation>0</Operation><Orientation>0</Orientation><Width WidthComput="0" WidthUnit="1" WidthSrc="1" WidthType="0">100</Width><Height HeightComput="0" HeightUnit="1" HeightSrc="1" HeightType="1">100</Height><ConstrainProportions>True</ConstrainProportions><HorizontalJustification>2</HorizontalJustification><VerticalJustification>2</VerticalJustification><HorizontalOffset HorizontalOffsetUnit="0" HorizontalOffsetDir="0">0</HorizontalOffset><VerticalOffset VerticalOffsetUnit="0" VerticalOffsetDir="0">0</VerticalOffset></Task><Task type="DeleteTagTask" enabled="True"><DelType>0</DelType><DelSpecTag>1</DelSpecTag></Task><Task type="SetTagTask" enabled="True"><TagType>58</TagType><IPTC_Keywords><![CDATA[a,b,c,d]]></IPTC_Keywords></Task><Task type="SaveAsTask" enabled="True"><FileName><![CDATA[<Original Name (Without Extension)>]]></FileName><PreserveStruct>False</PreserveStruct><CommonFolder><![CDATA[]]></CommonFolder><FileType></FileType><FilePath><![CDATA[<Source Folder>out]]></FilePath><FileExists>3</FileExists><DefaultOptions>True</DefaultOptions><BMPCompression>0</BMPCompression><BMPVersion>1</BMPVersion><JPEGColorSpace>2</JPEGColorSpace><JPEGDCTMethod>0</JPEGDCTMethod><JPEGCromaSubsampling>1</JPEGCromaSubsampling><JPEGOptimalHuffman>False</JPEGOptimalHuffman><JPEGQuality>85</JPEGQuality><PNGCompression>5</PNGCompression><PNGFilter>1</PNGFilter><PNGInterlaced>False</PNGInterlaced><J2000ColorSpace>1</J2000ColorSpace><J2000Rate>0/500</J2000Rate><PCXCompression>1</PCXCompression><HDPLossless>False</HDPLossless><HDPImageQuality>0/900</HDPImageQuality><TGACompressed>False</TGACompressed></Task></TaskList></Batch>
